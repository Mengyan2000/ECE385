    Mac OS X            	   2   |      �                                      ATTR       �   �                     �     com.apple.quarantine q/0082;63165632;Mail; 